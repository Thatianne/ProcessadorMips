library verilog;
use verilog.vl_types.all;
entity MemInstruction_TB is
end MemInstruction_TB;
