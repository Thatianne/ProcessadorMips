module Processor(clock)

IF IF ()

endmodule